library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity SPIhandler is
    port (
        clk : in std_logic;
        rst : in std_logic;
        sig
    );
end SPIhandler;

architecture rtl of SPIhandler is

begin

end architecture;